module top;
   test tb();
endmodule
