package payload_pkg;
   
class payload;
   bit [63:0] payload;
endclass

endpackage
