package PacketBad_pkg;
   import Packet_pkg;
class PacketBad extends Packet;
endclass
endpackage
