package Packet_bad_pkg;
   import Packet_pkg;
class Packet_bad extends Packet;
endclass
endpackage
